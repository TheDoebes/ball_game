

architecture behavior of game is
--signals

	signal ballx : integer := 0;
	signal bally : integer := 0;
	signal 

begin

--start with score logic

score:process(ballx, bally)